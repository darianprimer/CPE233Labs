`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Cal Poly SLO CPE 233
// Engineer: Darian Primer
// 
// Create Date: 02/05/2019 11:03:55 PM
// Description: RAT MCU
//////////////////////////////////////////////////////////////////////////////////


module RAT_MCU(
	input INTERUPT_IN, RESET, CLK,
	input [7:0] IN_PORT,
	output logic IO_STRB,
	output logic [7:0] OUT_PORT, PORT_ID
    );
	
	//OUTPUT FROM INTERUPT TO CONTROL UNIT
	logic I_OUT, INTERUPT_S;
	//OUTPUTS FROM CONTROL UNIT TO OTHER MODULES
	logic PC_LD_S, PC_INC_S, ALU_OPY_SEL_S, RF_WR_S, FLG_C_SET_S, FLG_C_CLR_S, FLG_C_LD_S, FLG_Z_LD_S, 
			RST_S, SP_LD_S, SP_INCR_S, SP_DECR_S, SCR_WE_S, SCR_DATA_SEL_S, I_SET_S, I_CLR_S, 
			FLG_LD_SEL_S, FLG_SHAD_LD_S;
	logic [1:0] PC_MUX_SEL_S, RF_WR_SEL_S, SCR_ADDR_SEL_S;
	logic [3:0] ALU_SEL_S;
	//OUTPUT FROM PROGRAM COUNTER TO OTHER MODULES
    logic [9:0] PC_COUNT_S;
	//OUTPUT FROM PROG_ROM TO OTHER MODULES
	logic [17:0] INSTRUCTION;
	//OUTPUT FROM REGISTER FILE TO OTHER MODULES
	logic [7:0] DX_OUT_S, DY_OUT_S;
	//OUTPUT FROM MUX FOR DIN OF REGISTER FILE
	logic [7:0] DIN_S;
    //OUTPUT FROM ALU TO OTHER MODULES
	logic [7:0] RESULT_S;
	logic C_S, Z_S;
	//OUTPUT FROM MUX FOR B OF ALU
	logic [7:0] B_S;
	//OUTPUT FROM FLAGS TO OTHER MODULES
	logic C_FLAG_S, Z_FLAG_S;
	//OUTPUT FROM STACK POINTER TO OTHER MODULES
	logic [7:0] DATASP_OUT_S;
	logic [7:0] DATASP2_OUT_S;
	//OUTPUT FROM SCRATCH RAM MUX1 TO SCRATCH RAM
	logic [9:0] DATASCR_IN_S;
	//OUTPUT FROM SCRATCH RAM MUX2 TO SCRATCH RAM
	logic [7:0] SCR_ADDR_S;
	//OUTPUT FROM SCRATCH RAM TO OTHER MODULES
	logic [9:0] DATASCR_OUT_S;
	
	assign DATASP2_OUT_S=DATASP_OUT_S-1;
	
	INTERUPT INTERUPT(.CLK(CLK), .SET(I_SET_S), .CLR(I_CLR_S), .OUT(I_OUT));
	
	assign INTERUPT_S=INTERUPT_IN&I_OUT;
	
    ControlUnit ControlUnit_inst(.C(C_FLAG_S), .Z(Z_FLAG_S), .INTERUPT(INTERUPT_S), .RESET(RESET), .CLK(CLK),  //INPUTS
							.OPCODE_HI_5(INSTRUCTION[17:13]), .OPCODE_LO_2(INSTRUCTION[1:0]), 			//INPUTS
							.PC_LD(PC_LD_S), .PC_INC(PC_INC_S), .ALU_OPY_SEL(ALU_OPY_SEL_S), 			//OUTPUTS
							.RF_WR(RF_WR_S), .FLG_C_SET(FLG_C_SET_S), .FLG_C_CLR(FLG_C_CLR_S),			//OUTPUTS
							.FLG_C_LD(FLG_C_LD_S), .FLG_Z_LD(FLG_Z_LD_S), .FLG_LD_SEL(FLG_LD_SEL_S), 	//OUTPUTS
							.FLG_SHAD_LD(FLG_SHAD_LD_S), .RST(RST_S), .I_SET(I_SET_S), .I_CLR(I_CLR_S),	//OUTPUTS
							.IO_STRB(IO_STRB), .PC_MUX_SEL(PC_MUX_SEL_S),								//OUTPUTS
							.RF_WR_SEL(RF_WR_SEL_S), .ALU_SEL(ALU_SEL_S), .SP_LD(SP_LD_S), 				//OUTPUTS
							.SP_INCR(SP_INCR_S), .SP_DECR(SP_DECR_S), .SCR_WE(SCR_WE_S), 				//OUTPUTS
							.SCR_DATA_SEL(SCR_DATA_SEL_S), .SCR_ADDR_SEL(SCR_ADDR_SEL_S));				//OUTPUTS
							
							
	
	
	PC_with_Mux PC_with_Mux(.FROM_IMMED(INSTRUCTION[12:3]), .FROM_STACK(DATASCR_OUT_S), .PC_MUX_SEL(PC_MUX_SEL_S), .PC_LD(PC_LD_S),
							.PC_INC(PC_INC_S), .RST(RST_S), .CLK(CLK), .PC_COUNT(PC_COUNT_S));

	
	
	ProgRom ProgRom(.PROG_CLK(CLK), .PROG_ADDR(PC_COUNT_S), .PROG_IR(INSTRUCTION));
	
	
	
	//MUX FOR DIN OF REGISTER FILE
	MUX_4IN MUX_4IN_inst1(.A(RESULT_S), .B(DATASCR_OUT_S), .C(DATASP_OUT_S), .D(IN_PORT), .MUX_SEL(RF_WR_SEL_S), .OUT(DIN_S));
	
	Register_File Register_File(.DIN(DIN_S), .ADRX(INSTRUCTION[12:8]), .ADRY(INSTRUCTION[7:3]), .RF_WR(RF_WR_S), .clk(CLK),
								.DX_OUT(DX_OUT_S), .DY_OUT(DY_OUT_S));
								
	
	//MUX FOR B OF ALU
	MUX_4IN MUX_4IN_inst2(.A(DY_OUT_S), .B(INSTRUCTION[7:0]), .C(), .D(), .MUX_SEL({1'b0, ALU_OPY_SEL_S}), .OUT(B_S));
								
	ALU ALU(.SEL(ALU_SEL_S), .A(DX_OUT_S), .B(B_S), .CIN(C_FLAG_S), .RESULT(RESULT_S), .C(C_S), .Z(Z_S));
	
	
	FLAGS FLAGS(.FLG_C_SET(FLG_C_SET_S), .FLG_C_CLR(FLG_C_CLR_S), .FLG_C_LD(FLG_C_LD_S), .FLG_Z_LD(FLG_Z_LD_S),
				.FLG_LD_SEL(FLG_LD_SEL_S), .FLG_SHAD_LD(FLG_SHAD_LD_S), .CLK(CLK), .C(C_S), .Z(Z_S),
				.C_FLG(C_FLAG_S), .Z_FLG(Z_FLAG_S));
				
	StackPointer StackPointer(.RST(RST_S), .LD(SP_LD_S), .INCR(SP_INCR_S), .DECR(SP_DECR_S), .DATA(DX_OUT_S), .CLK(CLK), .OUT(DATASP_OUT_S));
	
	//MUX FOR DATA_IN OF SCR
	MUX_2IN MUX_2IN_inst1(.A(DX_OUT_S), .B(PC_COUNT_S), .MUX_SEL(SCR_DATA_SEL_S), .OUT(DATASCR_IN_S));
	
	//MUX FOR ADDR OF SCR
	MUX_4IN MUX_4IN_inst3(.A(DY_OUT_S), .B(INSTRUCTION), .C(DATASP_OUT_S), .D(DATASP2_OUT_S), .MUX_SEL(SCR_ADDR_SEL_S), .OUT(SCR_ADDR_S));
	
	Scratch_RAM Scratch_RAM(.DATA_IN(DATASCR_IN_S), .SCR_WE(SCR_WE_S), .SCR_ADDR(SCR_ADDR_S), .clk(CLK), .DATA_OUT(DATASCR_OUT_S));
				
	assign OUT_PORT=DX_OUT_S;
	assign PORT_ID=INSTRUCTION[7:0];
	
endmodule
